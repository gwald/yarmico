pBAV       �       @       �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             @@        ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            